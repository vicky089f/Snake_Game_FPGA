`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 20.11.2021 11:50:18
// Design Name: 
// Module Name: square
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SnakeTopModule(
    input clk,
    input reset,
    input W,
    input A,
    input S,
    input D,
    output reg vga_hsync,
    output reg vga_vsync,
    output reg [3:0] vga_r,
    output reg [3:0] vga_g,
    output reg [3:0] vga_b
    );
    
    wire Clk_25,locked, Clk_Deb, Clk_Snake;
    wire [9:0] sx,sy;
    wire hsync,vsync,de,key,keypress;
    wire [2:0] Dir;
    wire snake_draw, head_draw, collide, food_draw;
    wire [7:0] Score;
    wire clk2, clk3, clk5, clk10;
    
    assign key = W || A || S || D || collide;
    Snake_Clocks snclk(clk, reset, clk2, clk3, clk5, clk10);
    
    clk_wiz_0 M1(.reset(reset), .clk_in(clk), .clk_out(Clk_25), .locked(locked));
    ClkDiv M2(clk, reset, Clk_Deb, Clk_Snake);
    debounce M3(Clk_Deb, reset, key, keypress);
    SnakeFSM M4(keypress, reset, W,A,S,D, collide, Dir);
    SnakeBody M5(/*Clk_Snake,*/ clk2, clk3, clk5, clk10, reset, sx, sy, Dir, head_draw, snake_draw, collide, food_draw, Score);
    VGA_480p M6(Clk_25, !locked, sx, sy, hsync, vsync, de);
    vio_0 M7(clk, Score);
    
    always@(posedge Clk_25)
    begin
        vga_hsync <= hsync;
        vga_vsync <= vsync;
        if(Dir != 5) begin
            vga_r <= !de ? 4'h0 : head_draw ? 4'hf : food_draw ? 4'hf : (snake_draw ? 4'h9 : 4'h2);
            vga_g <= !de ? 4'h0 : head_draw ? 4'ha : food_draw ? 4'h0 : (snake_draw ? 4'h9 : 4'h2);
            vga_b <= !de ? 4'h0 : head_draw ? 4'h6 : food_draw ? 4'h0 : (snake_draw ? 4'h9 : 4'h2);
        end
        else begin
            vga_r <= !de ? 4'h0 : 4'h0;
            vga_g <= !de ? 4'h0 : 4'h0;
            vga_b <= !de ? 4'h0 : 4'hf;
        end
    end
    
endmodule
